module sum (
  input wire [31:0] a, b, s
);
  assign s = a + b;
endmodule